`define MUX2