`define MUX1