`undef MUX1