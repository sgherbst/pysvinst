`undef MUX2