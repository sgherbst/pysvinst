module A;
endmodule