module A(
    b.in c
);
endmodule
